.subckt d g s pmos gm = 'gm' rds = 'rds' cgs = 'cgs'

gm d s s g gm
rds d s rds
cgs g s cgs

.ends pmos 

.ends